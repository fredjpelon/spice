A Berkeley SPICE3 compatible circuit
*
* This circuit contains only Berkeley SPICE3 components .
*
* The circuit is an AC coupled transistor amplifier with
* a sinewave input at node "1" , a gain of approximately -3.9 ,
* and output on node " coll ".
*
*.tran 1e-5 2e-3
*
vcc vcc 0 12.0
*vin 1 0 0.0 ac 1.0 sin (0 1 1k)
vin 1 0 0.0 ac 1.0 sin (0 1 2k)
ccouple 1 base 10uF
rbias1 vcc base 100k
rbias2 base 0 24k
q1 coll base emit generic
rcollector vcc coll 3.9k
remitter emit 0 1k
*
.model generic npn
*
.control
*tran 1e-5 2e-3
tran 1e-6 2e-3
set filetype=ascii
write npnout.txt v(base) v(coll)
.endc
.end